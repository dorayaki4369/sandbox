module Lesson1(switch, led);
	input switch;
	output led;
	
	assign led=switch;
endmodule